`timescale 1ns/1ps
//`include "alu.v"

module test();

reg[31:0] instruction;
reg[31:0] regA;
reg[31:0] regB;
wire[31:0] result;
wire[2:0] flags;

initial
begin
    $dumpfile("test.vcd");
    $dumpvars;
end

initial
begin
    $monitor("instruction=32'b%b, regA=32'b%b, regB=32'b%b,result=32'b%b, flags=3'b%b",instruction,regA,regB,result,flags);
    instruction=32'b0;
    regA=32'b0;
    regB=32'b0;

    #100
    $display("\n Add test#1(normal add)");
    instruction=32'b000000_00000_00001_00000_00000_100000;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Add test#2(overflow add)");
    instruction=32'b000000_00000_00001_00000_00000_100000;
    regA=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_1001;

    #100
    $display("\n Addu test");
    instruction=32'b000000_00000_00001_00000_00000_100001;
    regA=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_1001;

    #100
    $display("\n Sub test#1(normal sub)");
    instruction=32'b000000_00000_00001_00000_00000_100010;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Sub test#2(overflow sub)");
    instruction=32'b000000_00000_00001_00000_00000_100010;
    regA=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    regB=32'b1111_1111_1111_1111_1111_1111_1111_1111;

    #100
    $display("\n Subu test");
    instruction=32'b000000_00000_00001_00000_00000_100001;
    regA=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    regB=32'b1111_1111_1111_1111_1111_1111_1111_1111;

    #100
    $display("\n And test");
    instruction=32'b000000_00000_00001_00000_00000_100100;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0011;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0101;

    #100
    $display("\n Nor test");
    instruction=32'b000000_00000_00001_00000_00000_100111;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0011;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0101;

    #100
    $display("\n Or test");
    instruction=32'b000000_00000_00001_00000_00000_100101;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0011;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0101;

    #100
    $display("\n Xor test");
    instruction=32'b000000_00000_00001_00000_00000_100110;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0011;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0101;

    #100
    $display("\n Slt test#1(negative)");
    instruction=32'b000000_00000_00001_00000_00000_101010;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Slt test#2(non-negative)");
    instruction=32'b000000_00000_00001_00000_00000_101010;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Sltu test#1(negative)");
    instruction=32'b000000_00000_00001_00000_00000_101011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Sltu test#2(non-negative)");
    instruction=32'b000000_00000_00001_00000_00000_101011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Sll test");
    instruction=32'b000000_00000_00001_00000_00001_000000;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Sllv test");
    instruction=32'b000000_00000_00001_00000_00000_000100;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Srl test");
    instruction=32'b000000_00000_00001_00000_00001_000010;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    
    #100
    $display("\n Srlv test");
    instruction=32'b000000_00000_00001_00000_00000_000110;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Sra test");
    instruction=32'b000000_00000_00001_00000_00001_000011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Srav test");
    instruction=32'b000000_00000_00001_00000_00000_000111;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Addi test#1(normal addi)");
    instruction=32'b001000_00000_00001_0000_0000_0000_0001;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    #100
    $display("\n Addi test#2(overflow addi)");
    instruction=32'b001000_00000_00001_0000_0000_0000_0001;
    regA=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Addiu test");
    instruction=32'b001001_00000_00001_0000_0000_0000_0001;
    regA=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Andi test");
    instruction=32'b001001_00000_00001_0000_0000_0000_0011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Beq test#1");
    instruction=32'b000100_00000_00001_0000_0000_0000_0001;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Beq test#2");
    instruction=32'b000100_00000_00001_0000_0000_0000_0001;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;   

    #100
    $display("\n Bne test#1");
    instruction=32'b000101_00000_00001_0000_0000_0000_0001;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Bne test#2");
    instruction=32'b000101_00000_00001_0000_0000_0000_0001;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    #100
    $display("\n Ori test");
    instruction=32'b001101_00000_00001_0000_0000_0000_0011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Xori test");
    instruction=32'b001110_00000_00001_0000_0000_0000_0011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Slti test#1(negative)");
    instruction=32'b001010_00000_00001_0000_0000_0000_0001;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0000;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    #100
    $display("\n Slti test#2(non-negative)");
    instruction=32'b001010_00000_00001_0000_0000_0000_0000;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    #100
    $display("\n Sltiu test#1(negative)");
    instruction=32'b001011_00000_00001_0000_0000_0001_0000;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    #100
    $display("\n Sltiu test#2(non-negative)");
    instruction=32'b001011_00000_00001_0000_0000_0001_0000;
    regA=32'b0000_0000_0000_0000_0000_0000_1000_0000;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    #100
    $display("\n Lw test");
    instruction=32'b100011_00000_00001_0000_0000_0000_0011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $display("\n Sw test");
    instruction=32'b101011_00000_00001_0000_0000_0000_0011;
    regA=32'b0000_0000_0000_0000_0000_0000_0000_0101;
    regB=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    #100
    $stop;
end

alu u_add(
    .instruction(instruction),
    .regA(regA),
    .regB(regB),
    .result(result),
    .flags(flags)
);

endmodule